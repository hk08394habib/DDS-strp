// Copyright 2023 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.



module counter (input clk,
                input reset,
                output reg [3:0] count_out = 4'b1);

   always @(posedge clk) begin
      count_out <= count_out + 4'b1;
   end

   always @(negedge reset) begin
      count_out <= 4'b0;
   end


endmodule



